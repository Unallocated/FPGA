library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.uas.ALL;

entity text_bitmap is
	 Generic ( 
				red_width   : positive := 3;
				green_width : positive := 3;
				blue_width  : positive := 2
				);
    Port ( 
	      clk   : in  STD_LOGIC;
         rst   : in  STD_LOGIC;
         hs    : out  STD_LOGIC;
         vs    : out  STD_LOGIC;
         red   : out  STD_LOGIC_VECTOR (red_width-1 downto 0);
         green : out  STD_LOGIC_VECTOR (green_width-1 downto 0);
         blue  : out  STD_LOGIC_VECTOR (blue_width-1 downto 0)
			);
end text_bitmap;

architecture Behavioral of text_bitmap is

	COMPONENT vga_configurable
	Generic ( 
			  config      : vga_timing;
			  red_width   : positive;
			  green_width : positive;
			  blue_width  : positive
			  );
	PORT(
		clk      : IN std_logic;
		rst      : IN std_logic;
		blue_in  : IN std_logic_vector;
		red_in   : IN std_logic_vector;
		green_in : IN std_logic_vector;          
		hs       : OUT std_logic;
		vs       : OUT std_logic;
		green    : OUT std_logic_vector;
		red      : OUT std_logic_vector;
		blue     : OUT std_logic_vector;
		x_pos    : OUT integer range -1 to config.horizontal_video - 1;
		y_pos    : OUT integer range -1 to config.vertical_video - 1
		);
	END COMPONENT;
	
	-- Nexys3
--	COMPONENT nexys3_clock
--	PORT(
--	  CLK_IN1  : in  std_logic;
--	  CLK_OUT1 : out std_logic
--	    );
--	END COMPONENT;
	
	-- Mojo
	COMPONENT mojo_clock
	PORT(
	  CLK_IN1  : in  std_logic;
	  CLK_OUT1 : out std_logic
	    );
	END COMPONENT;
	
	-- Basys2
--	COMPONENT clock
--	PORT(
--		CLKIN_IN        : IN std_logic;          
--		CLKFX_OUT       : OUT std_logic;
--		CLKIN_IBUFG_OUT : OUT std_logic;
--		CLK0_OUT        : OUT std_logic
--		 );
--	END COMPONENT;
	
	constant vga_config : vga_timing := vga_25mhz_640x480;
	
	signal vga_clk : std_logic;
	
	signal red_buf   : std_logic_vector(red_width - 1 downto 0)   := (others => '1');
	signal green_buf : std_logic_vector(green_width - 1 downto 0) := (others => '0');
	signal blue_buf  : std_logic_vector(blue_width - 1 downto 0)  := (others => '0');
	
	signal x_pos : integer range -1 to vga_config.horizontal_video - 1;
	signal y_pos : integer range -1 to vga_config.vertical_video - 1;
	
	
	type bitmap_type is array (0 to 19) of std_logic_vector(0 to 199);
	constant bitmap : bitmap_type := 
	(
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
		("00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000110011000"),
		("01111111010000000100000000000001000000000000000000000000010000000000000000000100000000000000001000000000000000000000000000010000000100100000000000000000000000000000000000000000010000000000001000100000"),
		("00001000010000000000000000000000000000000000000000000000010000000000000000000100000000000000001000000000000000000000000000010000000000100000000000000000000000000000000000000000010000000000001000100000"),
		("00001000010111000100011100000001000111000000001111000000111100011110000111001111000000011110011110000011110111001000010000011111000101111001111011100001111000111110000000011100111100100001011111111000"),
		("00001000011000100100100010000001001000100000010000100000010000110011001000100100000000110011001000000010001000101000010000011001100100100001000100010010000100110011000000100010010000100001001000100000"),
		("00001000010000100100100000000001001000000000000000100000010000100001001000000100000000100001001000000010001000100100100000010000100100100001000100010000000100100001000000100000010000100001001000100000"),
		("00001000010000100100011100000001000111000000001111100000010000111111000111000100000000100001001000000010001000100100100000010000100100100001000100010001111100100001000000011100010000100001001000100000"),
		("00001000010000100100000010000001000000100000010000100000010000100000000000100100000000100001001000000010001000100010100000010000100100100001000100010010000100100001000000000010010000100001001000100000"),
		("00001000010000100100100010000001001000100000010001100000010000110001001000100100000000110011001000000010001000100011000000011001100100100001000100010010001100110011000000100010010000100011001000100000"),
		("00001000010000100100011100000001000111000000001110100000011100011110000111000111000000011110001000000010001000100001000000011111000100111001000100010001110100111110000000011100011100011101001000100000"),
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000"),
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000"),
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000100000000000000000000000000000000000000000"),
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
		("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111")
	);

begin

	process(vga_clk)
	begin
		if(rising_edge(vga_clk)) then
			if(x_pos - 100 > -1 and y_pos - 100 > -1 and x_pos - 100 < bitmap(0)'high + 1
					and y_pos - 100 < bitmap'high + 1) then
				if(bitmap(y_pos - 100)(x_pos - 100) = '1') then
					red_buf <= (others => '1');
				else
					red_buf <= (others => '0');
				end if;
			else
				red_buf <= (others => '0');
			end if;
		end if;
	end process;

	-- Nexys3
--	Inst_clock : nexys3_clock PORT MAP(
--		CLK_IN1 => clk,
--		CLK_OUT1 => vga_clk
--	);
	
	-- Mojo
	Inst_clock : mojo_clock PORT MAP(
		CLK_IN1 => clk,
		CLK_OUT1 => vga_clk
	);
	
	-- Basys2
--	Inst_clock: clock PORT MAP(
--		CLKIN_IN        => clk,
--		CLKFX_OUT       => vga_clk,
--		CLKIN_IBUFG_OUT => open,
--		CLK0_OUT        => open
--	);

	Inst_vga_configurable: vga_configurable 
	GENERIC MAP(
		config      => vga_25mhz_640x480,
		red_width   => red_width,
		green_width => green_width,
		blue_width  => blue_width
	)
	PORT MAP(
		clk      => vga_clk,
		rst      => rst,
		hs       => hs,
		vs       => vs,
		green    => green,
		red      => red,
		blue     => blue,
		x_pos    => x_pos,
		y_pos    => y_pos,
		blue_in  => blue_buf,
		red_in   => red_buf,
		green_in => green_buf
	);

end Behavioral;

